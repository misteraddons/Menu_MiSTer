//============================================================================
//
//  Menu for MiSTer.
//  Copyright (C) 2017-2020 Sorgelig
//
//
//  This program is free software; you can redistribute it and/or modify it
//  under the terms of the GNU General Public License as published by the Free
//  Software Foundation; either version 2 of the License, or (at your option)
//  any later version.
//
//  This program is distributed in the hope that it will be useful, but WITHOUT
//  ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
//  FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License for
//  more details.
//
//  You should have received a copy of the GNU General Public License along
//  with this program; if not, write to the Free Software Foundation, Inc.,
//  51 Franklin Street, Fifth Floor, Boston, MA 02110-1301 USA.
//
//============================================================================

module emu
(
	//Master input clock
	input         CLK_50M,

	//Async reset from top-level module.
	//Can be used as initial reset.
	input         RESET,

	//Must be passed to hps_io module
	inout  [48:0] HPS_BUS,

	//Base video clock. Usually equals to CLK_SYS.
	output        CLK_VIDEO,

	//Multiple resolutions are supported using different CE_PIXEL rates.
	//Must be based on CLK_VIDEO
	output        CE_PIXEL,

	//Video aspect ratio for HDMI. Most retro systems have ratio 4:3.
	//if VIDEO_ARX[12] or VIDEO_ARY[12] is set then [11:0] contains scaled size instead of aspect ratio.
	output [12:0] VIDEO_ARX,
	output [12:0] VIDEO_ARY,

	output  [7:0] VGA_R,
	output  [7:0] VGA_G,
	output  [7:0] VGA_B,
	output        VGA_HS,
	output        VGA_VS,
	output        VGA_DE,    // = ~(VBlank | HBlank)
	output        VGA_F1,
	output [1:0]  VGA_SL,
	output        VGA_SCALER, // Force VGA scaler
	output        VGA_DISABLE, // analog out is off

	input  [11:0] HDMI_WIDTH,
	input  [11:0] HDMI_HEIGHT,
	output        HDMI_FREEZE,
	output        HDMI_BLACKOUT,

`ifdef MISTER_FB
	// Use framebuffer in DDRAM
	// FB_FORMAT:
	//    [2:0] : 011=8bpp(palette) 100=16bpp 101=24bpp 110=32bpp
	//    [3]   : 0=16bits 565 1=16bits 1555
	//    [4]   : 0=RGB  1=BGR (for 16/24/32 modes)
	//
	// FB_STRIDE either 0 (rounded to 256 bytes) or multiple of pixel size (in bytes)
	output        FB_EN,
	output  [4:0] FB_FORMAT,
	output [11:0] FB_WIDTH,
	output [11:0] FB_HEIGHT,
	output [31:0] FB_BASE,
	output [13:0] FB_STRIDE,
	input         FB_VBL,
	input         FB_LL,
	output        FB_FORCE_BLANK,

`ifdef MISTER_FB_PALETTE
	// Palette control for 8bit modes.
	// Ignored for other video modes.
	output        FB_PAL_CLK,
	output  [7:0] FB_PAL_ADDR,
	output [23:0] FB_PAL_DOUT,
	input  [23:0] FB_PAL_DIN,
	output        FB_PAL_WR,
`endif
`endif

	output        LED_USER,  // 1 - ON, 0 - OFF.

	// b[1]: 0 - LED status is system status OR'd with b[0]
	//       1 - LED status is controled solely by b[0]
	// hint: supply 2'b00 to let the system control the LED.
	output  [1:0] LED_POWER,
	output  [1:0] LED_DISK,

	// I/O board button press simulation (active high)
	// b[1]: user button
	// b[0]: osd button
	output  [1:0] BUTTONS,

	input         CLK_AUDIO, // 24.576 MHz
	output [15:0] AUDIO_L,
	output [15:0] AUDIO_R,
	output        AUDIO_S,   // 1 - signed audio samples, 0 - unsigned
	output  [1:0] AUDIO_MIX, // 0 - no mix, 1 - 25%, 2 - 50%, 3 - 100% (mono)

	//ADC
	inout   [3:0] ADC_BUS,

	//SD-SPI
	output        SD_SCK,
	output        SD_MOSI,
	input         SD_MISO,
	output        SD_CS,
	input         SD_CD,

	//High latency DDR3 RAM interface
	//Use for non-critical time purposes
	output        DDRAM_CLK,
	input         DDRAM_BUSY,
	output  [7:0] DDRAM_BURSTCNT,
	output [28:0] DDRAM_ADDR,
	input  [63:0] DDRAM_DOUT,
	input         DDRAM_DOUT_READY,
	output        DDRAM_RD,
	output [63:0] DDRAM_DIN,
	output  [7:0] DDRAM_BE,
	output        DDRAM_WE,

	//SDRAM interface with lower latency
	output        SDRAM_CLK,
	output        SDRAM_CKE,
	output [12:0] SDRAM_A,
	output  [1:0] SDRAM_BA,
	inout  [15:0] SDRAM_DQ,
	output        SDRAM_DQML,
	output        SDRAM_DQMH,
	output        SDRAM_nCS,
	output        SDRAM_nCAS,
	output        SDRAM_nRAS,
	output        SDRAM_nWE,

`ifdef MISTER_DUAL_SDRAM
	//Secondary SDRAM
	//Set all output SDRAM_* signals to Z ASAP if SDRAM2_EN is 0
	input         SDRAM2_EN,
	output        SDRAM2_CLK,
	output [12:0] SDRAM2_A,
	output  [1:0] SDRAM2_BA,
	inout  [15:0] SDRAM2_DQ,
	output        SDRAM2_nCS,
	output        SDRAM2_nCAS,
	output        SDRAM2_nRAS,
	output        SDRAM2_nWE,
`endif

	input         UART_CTS,
	output        UART_RTS,
	input         UART_RXD,
	output        UART_TXD,
	output        UART_DTR,
	input         UART_DSR,

	// Open-drain User port.
	// 0 - D+/RX
	// 1 - D-/TX
	// 2..6 - USR2..USR6
	// Set USER_OUT to 1 to read from USER_IN.
	input   [6:0] USER_IN,
	output  [6:0] USER_OUT,

	input         OSD_STATUS
);

assign ADC_BUS  = 'Z;
assign {UART_RTS, UART_DTR} = 0;
assign {SD_SCK, SD_MOSI, SD_CS} = 'Z;

assign DDRAM_CLK = clk_sys;
assign CE_PIXEL  = ce_pix;

assign VGA_SL = 0;
assign VGA_F1 = 0;
assign VIDEO_ARX = 0;
assign VIDEO_ARY = 0;
assign VGA_SCALER= 0;
assign VGA_DISABLE = 0;

assign AUDIO_MIX = 0;
assign HDMI_FREEZE = 0;
assign HDMI_BLACKOUT = 0;

assign LED_DISK = 0;
assign LED_POWER[1]= 1;
assign BUTTONS = 0;

reg  [26:0] act_cnt;
always @(posedge clk_sys) act_cnt <= act_cnt + 1'd1; 
assign LED_USER    = FB ? led[0] : act_cnt[26]  ? act_cnt[25:18]  > act_cnt[7:0]  : act_cnt[25:18]  <= act_cnt[7:0];

wire [26:0] act_cnt2 = {~act_cnt[26],act_cnt[25:0]};
assign LED_POWER[0]= FB ? led[2] : act_cnt2[26] ? act_cnt2[25:18] > act_cnt2[7:0] : act_cnt2[25:18] <= act_cnt2[7:0];


`include "build_id.v" 
localparam CONF_STR = {
	"MENU;UART31250,MIDI;",
	"-;",
	"T0,Show CFG Debug;",
	"-;", 
	"V,v",`BUILD_DATE 
};

wire forced_scandoubler;
wire [31:0] status;

hps_io #(.CONF_STR(CONF_STR)) hps_io
(
	.clk_sys(clk_sys),
	.HPS_BUS(HPS_BUS),
	.forced_scandoubler(forced_scandoubler),
	.status(status),
	.status_menumask(cfg)
);

////////////////////   CLOCKS   ///////////////////
wire locked, clk_sys;
pll pll
(
	.refclk(CLK_50M),
	.rst(0),
	.outclk_0(clk_sys),
	.outclk_1(CLK_VIDEO),
	.locked(locked)
);


/////////////////////   SDRAM   ///////////////////
//
// Helper functionality:
//    SDRAM and DDR3 RAM are being cleared while this core is working.
//    some cores behave incorrectly if started with non-clean RAM.

sdram sdr
(
	.*,
	.init(~locked),
	.clk(clk_sys),
	.addr(sdram_addr),
	.wtbt(3),
	.dout(sdram_dout),
	.din(sdram_din),
	.rd(sdram_rd),
	.we(sdram_we),
	.ready(sdram_ready)
);

reg  [26:0] sdram_addr;
wire        sdram_ready;
wire [15:0] sdram_dout;
reg  [15:0] sdram_din;
reg         sdram_we;
reg         sdram_rd;

`ifdef MISTER_DUAL_SDRAM
// Secondary SDRAM interface for capacity testing
reg  [26:0] sdram2_addr;
wire        sdram2_ready;
wire [15:0] sdram2_dout;
reg  [15:0] sdram2_din;
reg         sdram2_we;
reg         sdram2_rd;
`endif

reg  [15:0] cfg = 0;

always @(posedge clk_sys) begin
	reg [5:0] state = 0;

	sdram_rd <= 0;
	sdram_we <= 0;
`ifdef MISTER_DUAL_SDRAM
	sdram2_rd <= 0;
	sdram2_we <= 0;
`endif

	if(RESET) begin
		state <= 0;
		cfg <= 0;  // All configuration bits start at 0
	end
	else begin
		case(state)
			// Primary SDRAM testing (states 0-15)
			0: if(sdram_ready) begin
					cfg <= 0;  // Clear all configuration bits
					state      <= state+1'd1;
				end
			1: begin
					sdram_addr <= 'h4000000;
					sdram_din  <= 3128;
					sdram_we   <= 1;
					state      <= state+1'd1;
				end
			2: state <= state+1'd1;
			3: if(sdram_ready) begin
					sdram_addr <= 'h2000000;
					sdram_din  <= 2064;
					sdram_we   <= 1;
					state      <= state+1'd1;
				end
			4: state <= state+1'd1;
			5: if(sdram_ready) begin
					sdram_addr <= 'h0000000;
					sdram_din  <= 1032;
					sdram_we   <= 1;
					state      <= state+1'd1;
				end
			6: state <= state+1'd1;
			7: if(sdram_ready) begin
					sdram_addr <= 'h1000000;
					sdram_din  <= 12345;
					sdram_we   <= 1;
					state      <= state+1'd1;
				end
			8: state <= state+1'd1;
			9: if(sdram_ready) begin
					sdram_addr <= 'h4000000;
					sdram_rd   <= 1;
					state      <= state+1'd1;
				end
			10: state <= state+1'd1;
			11: if(sdram_ready) begin
					cfg[2]     <= (sdram_dout == 3128);
					sdram_addr <= 'h2000000;
					sdram_rd   <= 1;
					state      <= state+1'd1;
				end
			12: state <= state+1'd1;
			13: if(sdram_ready) begin
					cfg[1]     <= (sdram_dout == 2064);
					sdram_addr <= 'h0000000;
					sdram_rd   <= 1;
					state      <= state+1'd1;
				end
			14: state <= state+1'd1;
			15: if(sdram_ready) begin
					cfg[0]     <= (sdram_dout == 1032);
					//cfg[15] <= 1;  // Primary SDRAM present flag
					state      <= state+1'd1;
				end

`ifdef MISTER_DUAL_SDRAM
			// Secondary SDRAM testing (states 16-31)
			//16: if(sdram_ready) begin
			//		cfg <= 0;  // Clear all configuration bits
			//		state      <= state+1'd1;
			//	end
			
			//16: if(SDRAM2_EN && sdram2_ready) begin
			/*
			16: begin
					//cfg[7] <= 1;  // Debug: mark that we reached state 16
					if(sdram2_ready) begin
						// Hardware presence test - write distinctive pattern  
						sdram2_addr <= 'h0800000;  // Use address 8MB for presence test
						sdram2_din  <= 16'hA5A5;   // Distinctive test pattern
						sdram2_we   <= 1;
						cfg[5:3]    <= 3'd0;       // Clear secondary bits
						state       <= state+1'd1;
					end
					else begin
						// No secondary SDRAM hardware, skip to completion  
						cfg[6:3]   <= 4'd0;  // Clear secondary bits and presence flag
						cfg[15]    <= 1;
						state      <= state+16;
					end
				end
				*/
			16: if(sdram2_ready) begin
					sdram2_addr <= 'h4000000;
					sdram2_din  <= 3128;
					sdram2_we   <= 1;
					state      <= state+1'd1;
				end
			17: state <= state+1'd1;
			18: if(sdram2_ready) begin
					sdram2_addr <= 'h2000000;
					sdram2_din  <= 2064;
					sdram2_we   <= 1;
					state      <= state+1'd1;
				end
			19: state <= state+1'd1;
			20: if(sdram2_ready) begin
					sdram2_addr <= 'h0000000;
					sdram2_din  <= 1032;
					sdram2_we   <= 1;
					state      <= state+1'd1;
				end
			21: state <= state+1'd1;
			22: if(sdram2_ready) begin
					sdram2_addr <= 'h1000000;
					sdram2_din  <= 12345;
					sdram2_we   <= 1;
					state      <= state+1'd1;
				end
			23: state <= state+1'd1;
			24: if(sdram2_ready) begin
					sdram2_addr <= 'h4000000;
					sdram2_rd   <= 1;
					state      <= state+1'd1;
				end
			25: state <= state+1'd1;
			26: if(sdram2_ready) begin
					cfg[5]     <= (sdram2_dout == 3128);
					sdram2_addr <= 'h2000000;
					sdram2_rd   <= 1;
					cfg[6]   <= 1;    // Hardware present flag
					state      <= state+1'd1;
				end
			27: state <= state+1'd1;
			28: if(sdram2_ready) begin
					cfg[4]     <= (sdram2_dout == 2064);
					sdram2_addr <= 'h0000000;
					sdram2_rd   <= 1;
					cfg[6]   <= 1;    // Hardware present flag
					state      <= state+1'd1;
				end
			29: state <= state+1'd1;
			30: if(sdram2_ready) begin
					cfg[3]     <= (sdram2_dout == 1032);
					cfg[6]   <= 1;    // Secondary SDRAM present flag
					state      <= state+1'd1;
				end
`endif
			31: begin
					cfg[15] <= 1;     // Primary SDRAM present flag or test complete?
					sdram_addr <= addr[24:0];
					sdram_din  <= 0;
					sdram_we   <= we;
					sdram2_addr <= addr[24:0];
					sdram2_din  <= 0;
					sdram2_we   <= we;
				end

/*
			16: if(SDRAM2_EN && sdram2_ready) begin
					// Hardware presence test - write distinctive pattern  
					sdram2_addr <= 'h0800000;  // Use address 8MB for presence test
					sdram2_din  <= 16'hA5A5;   // Distinctive test pattern
					sdram2_we   <= 1;
					cfg[5:3]    <= 3'd0;       // Clear secondary bits
					state       <= state+1'd1;
				end
				else begin
					// No secondary SDRAM hardware, skip to completion  
					cfg[6:3]   <= 4'd0;  // Clear secondary bits and presence flag
					cfg[15]    <= 1;
					state      <= state+16;
				end
			17: state <= state+1'd1;
			18: if(sdram2_ready) begin
					// Read back the presence test pattern
					sdram2_addr <= 'h0800000;  // Read from presence test address
					sdram2_rd   <= 1;
					state      <= state+1'd1;
				end
			19: state <= state+1'd1;
			20: if(sdram2_ready) begin
					// Verify hardware presence before capacity testing
					if (sdram2_dout == 16'hA5A5) begin
						// Hardware present, start capacity testing with safe boundary
						sdram2_addr <= 'h4000000;  // 64MB boundary (same as primary)
						sdram2_din  <= 3128;       // Same pattern as primary
						sdram2_we   <= 1;
						state      <= state+1'd1;
					end
					else begin
						// Hardware not present - skip testing
						cfg[6:3] <= 4'd0;  // Clear secondary bits and presence flag
						cfg[15]  <= 1;
						state    <= state+12;
					end
				end
			21: state <= state+1'd1;
			22: if(sdram2_ready) begin
					sdram2_addr <= 'h2000000;  // 32MB boundary (same as primary)
					sdram2_din  <= 2064;       // Same pattern as primary
					sdram2_we   <= 1;
					state      <= state+1'd1;
				end
			23: state <= state+1'd1;
			24: if(sdram2_ready) begin
					sdram2_addr <= 'h0000000;  // Base address (same as primary)
					sdram2_din  <= 1032;       // Same pattern as primary  
					sdram2_we   <= 1;
					state      <= state+1'd1;
				end
			25: state <= state+1'd1;
			26: if(sdram2_ready) begin
					sdram2_addr <= 'h4000000;  // Read from 64MB boundary (same as primary)
					sdram2_rd   <= 1;
					state      <= state+1'd1;
				end
			27: state <= state+1'd1;
			28: if(sdram2_ready) begin
					cfg[5]      <= (sdram2_dout == 3128);  // 64MB+ test (same as primary cfg[2])
					sdram2_addr <= 'h2000000;  // Read from 32MB boundary (same as primary)
					sdram2_rd   <= 1;
					state      <= state+1'd1;
				end
			29: state <= state+1'd1;
			30: if(sdram2_ready) begin
					cfg[4]      <= (sdram2_dout == 2064);  // 32MB+ test (same as primary cfg[1])
					sdram2_addr <= 'h0000000;  // Read from base address (same as primary)
					sdram2_rd   <= 1;
					state      <= state+1'd1;
				end
			31: if(sdram2_ready) begin
					cfg[3]      <= (sdram2_dout == 1032);  // Base test (same as primary cfg[0])
					// Final secondary SDRAM validation and encoding
					// Now we have: cfg[5]=64MB+, cfg[4]=32MB+, cfg[3]=base
					if (cfg[5] && cfg[4] && (sdram2_dout == 1032)) begin
						// All tests passed = 128MB
						cfg[5:3] <= 3'd7; // 111 = 128MB
						cfg[6]   <= 1;    // Hardware present flag
					end
					else if (cfg[5] && cfg[4]) begin
						// 64MB+ and 32MB+ tests passed = 64MB
						cfg[5:3] <= 3'd3; // 011 = 64MB
						cfg[6]   <= 1;    // Hardware present flag
					end
					else if (cfg[4]) begin
						// Only 32MB+ test passed = 32MB
						cfg[5:3] <= 3'd1; // 001 = 32MB
						cfg[6]   <= 1;    // Hardware present flag
					end
					else begin
						// No tests passed = no hardware
						cfg[5:3] <= 3'd0; // 000 = no SDRAM
						cfg[6]   <= 0;    // No hardware present
					end
					cfg[15]     <= 1;  // Test complete
					state       <= state+1'd1;
				end
`else
			16: begin
					cfg[15]    <= 1;
					state      <= state+1'd1;
				end
`endif
			32: begin
					sdram_addr <= addr[24:0];
					sdram_din  <= 0;
					sdram_we   <= we;
				end
*/
		endcase
	end
end

ddram ddr
(
	.*,
	.reset(RESET),
   .dout(),
   .din(0),
   .rd(0),
   .ready()
);

`ifdef MISTER_DUAL_SDRAM
// Secondary SDRAM controller for capacity testing
sdram sdram2
(
	.init(~locked),
	.clk(clk_sys),
	.addr(sdram2_addr),
	.wtbt(3),
	.dout(sdram2_dout),
	.din(sdram2_din),
	.rd(sdram2_rd),
	.we(sdram2_we),
	.ready(sdram2_ready),

	// Secondary SDRAM pins  
	.SDRAM_DQ(SDRAM2_DQ),
	.SDRAM_A(SDRAM2_A),
	.SDRAM_BA(SDRAM2_BA),
	.SDRAM_nCS(SDRAM2_nCS),
	.SDRAM_nWE(SDRAM2_nWE),
	.SDRAM_nRAS(SDRAM2_nRAS),
	.SDRAM_nCAS(SDRAM2_nCAS),
	.SDRAM_CLK(SDRAM2_CLK),
	.SDRAM_CKE(),  // Not connected for secondary
	.SDRAM_DQML(), // Not connected for secondary  
	.SDRAM_DQMH()  // Not connected for secondary
);
`endif

reg        we;
reg [28:0] addr = 0;

always @(posedge clk_sys) begin
	reg [4:0] cnt = 9;

	if(~RESET & cfg[15]) begin
		cnt <= cnt + 1'b1;
		we <= &cnt;
		if(cnt == 8) addr <= addr + 1'd1;
	end
end

////////////////////////////  MT32pi  ////////////////////////////////// 

//
// Pin | USB Name | Signal
// ----+----------+--------------
// 0   | D+       | I/O I2C_SDA / RX (midi in)
// 1   | D-       | O   TX (midi out)
// 2   | TX-      | I   I2S_WS (1 == right)
// 3   | GND_d    | I   I2C_SCL
// 4   | RX+      | I   I2S_BCLK
// 5   | RX-      | I   I2S_DAT
// 6   | TX+      | -   none
//

reg [15:0] mt32_i2s_r, mt32_i2s_l;
wire midi_rx;

assign AUDIO_L = mt32_i2s_l;
assign AUDIO_R = mt32_i2s_r;
assign AUDIO_S = 1;

assign USER_OUT[0]   = 1;
assign USER_OUT[1]   = UART_RXD;
assign USER_OUT[6:2] = '1;
assign UART_TXD      = midi_rx;


//
// crossed/straight cable selection
//

generate
genvar i;
for(i = 0; i<2; i++) begin : clk_rate
	wire clk_in = i ? USER_IN[6] : USER_IN[4];
	reg [4:0] cnt;
	always @(posedge CLK_AUDIO) begin : clkr
		reg       clk_sr, clk, old_clk;
		reg [4:0] cnt_tmp;

		clk_sr <= clk_in;
		if (clk_sr == clk_in) clk <= clk_sr;

		if(~&cnt_tmp) cnt_tmp <= cnt_tmp + 1'd1;
		else cnt <= '1;

		old_clk <= clk;
		if(~old_clk & clk) begin
			cnt <= cnt_tmp;
			cnt_tmp <= 0;
		end
	end
end

reg crossed;
always @(posedge CLK_AUDIO) crossed <= (clk_rate[0].cnt <= clk_rate[1].cnt);
endgenerate

wire   i2s_ws   = crossed ? USER_IN[2] : USER_IN[5];
wire   i2s_data = crossed ? USER_IN[5] : USER_IN[2];
wire   i2s_bclk = crossed ? USER_IN[4] : USER_IN[6];
assign midi_rx  = crossed ? USER_IN[6] : USER_IN[4];

always @(posedge CLK_AUDIO) begin : i2s_proc
	reg [15:0] i2s_buf = 0;
	reg  [4:0] i2s_cnt = 0;
	reg        clk_sr;
	reg        i2s_clk = 0;
	reg        old_clk, old_ws;
	reg        i2s_next = 0;

	// Debounce clock
	clk_sr <= i2s_bclk;
	if (clk_sr == i2s_bclk) i2s_clk <= clk_sr;

	// Latch data and ws on rising edge
	old_clk <= i2s_clk;
	if (i2s_clk && ~old_clk) begin

		if (~i2s_cnt[4]) begin
			i2s_cnt <= i2s_cnt + 1'd1;
			i2s_buf[~i2s_cnt[3:0]] <= i2s_data;
		end

		// Word Select will change 1 clock before the new word starts
		old_ws <= i2s_ws;
		if (old_ws != i2s_ws) i2s_next <= 1;
	end

	if (i2s_next) begin
		i2s_next <= 0;
		i2s_cnt <= 0;
		i2s_buf <= 0;

		if (i2s_ws) mt32_i2s_l <= i2s_buf;
		else        mt32_i2s_r <= i2s_buf;
	end
	
	if (RESET) begin
		i2s_buf    <= 0;
		mt32_i2s_l <= 0;
		mt32_i2s_r <= 0;
	end
end

/////////////////////   VIDEO   ///////////////////

localparam lfsr_n = 63;

wire PAL = status[4];
wire FB  = status[5];
wire [2:0] led = status[8:6];

reg   [9:0] hc;
reg   [9:0] vc;
reg   [9:0] vvc;

reg  [lfsr_n:0] rnd_reg;
wire [lfsr_n:0] rnd;

wire  [5:0] rnd_c = {rnd_reg[0],rnd_reg[1],rnd_reg[2],rnd_reg[2],rnd_reg[2],rnd_reg[2]};

lfsr #(lfsr_n) random(rnd);

always @(posedge CLK_VIDEO) begin
	if(forced_scandoubler) ce_pix <= 1;
		else ce_pix <= ~ce_pix;

	if(ce_pix) begin
		if(hc == 637) begin
			hc <= 0;
			if(vc == (PAL ? (forced_scandoubler ? 623 : 311) : (forced_scandoubler ? 523 : 261))) begin 
				vc <= 0;
				vvc <= vvc + 9'd6;
			end else begin
				vc <= vc + 1'd1;
			end
		end else begin
			hc <= hc + 1'd1;
		end

		rnd_reg <= rnd;
	end
end

reg HBlank;
reg HSync;
reg VBlank;
reg VSync;

reg ce_pix;
always @(posedge CLK_VIDEO) begin
	if (hc == 529) HBlank <= 1;
		else if (hc == 0) HBlank <= 0;

	if (hc == 544) begin
		HSync <= 1;

		if(PAL) begin
			if(vc == (forced_scandoubler ? 609 : 304)) VSync <= 1;
				else if (vc == (forced_scandoubler ? 617 : 308)) VSync <= 0;

			if(vc == (forced_scandoubler ? 601 : 300)) VBlank <= 1;
				else if (vc == 0) VBlank <= 0;
		end
		else begin
			if(vc == (forced_scandoubler ? 490 : 245)) VSync <= 1;
				else if (vc == (forced_scandoubler ? 496 : 248)) VSync <= 0;

			if(vc == (forced_scandoubler ? 480 : 240)) VBlank <= 1;
				else if (vc == 0) VBlank <= 0;
		end
	end
	
	if (hc == 590) HSync <= 0;
end

reg  [7:0] cos_out;
wire [5:0] cos_g = cos_out[7:3]+6'd32;
cos cos(vvc + {vc>>forced_scandoubler, 2'b00}, cos_out);

wire [7:0] comp_v = (cos_g >= rnd_c) ? {cos_g - rnd_c, 2'b00} : 8'd0;

assign VGA_DE  = ~(HBlank | VBlank);
assign VGA_HS  = HSync;
assign VGA_VS  = VSync;
assign VGA_G   = comp_v;
assign VGA_R   = comp_v;
assign VGA_B   = comp_v;

endmodule
